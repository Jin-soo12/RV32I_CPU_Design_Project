`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];
    initial begin  //Simulation을 위한 임의의 명령어 할당
        $readmemh("code.mem", rom);
        /*
        //rom[x] = 32'b func7_rs2  _rs1  _f3 _rd   _op   // R-Type
        rom[0] =  32'b0000000_00010_00001_000_00011_0110011;// add x3, x1, x2 -> x3 = x1(-100) + x2(3)
        rom[1] =  32'b0100000_00010_00001_000_00100_0110011;// sub x4, x1, x2 -> x4 = x1(-100) - x2(3)
        rom[2] =  32'b0000000_00010_00001_001_00101_0110011;// sll x5, x1, x2 -> x5 = x1(-100) << x2(3)
        rom[3] =  32'b0000000_00010_00001_101_00110_0110011;// srl x6, x1, x2 -> x6 = x1(-100) >> x2(3)
        rom[4] =  32'b0100000_00010_00001_101_00111_0110011;// sra x7, x1, x2 -> x7 = x1(-100) >>> x2(3)
        rom[5] =  32'b0000000_00010_00001_010_01000_0110011;// slt x8, x1, x2 -> x8 = x1(-100) < x2(3) ? 1 : 0
        rom[6] =  32'b0000000_00010_00001_011_01001_0110011;// sltu x9, x1, x2 -> x9 = x1(-100) < x2(3) ? 1 : 0
        rom[7] =  32'b0000000_00010_00001_100_01010_0110011;// xor x10, x1, x2 -> x10 = x1(-100) ^ x2(3)
        rom[8] =  32'b0000000_00010_00001_110_01011_0110011;// or x11, x1, x2 -> x11 = x1(-100) | x2(3)
        rom[9] =  32'b0000000_00010_00001_111_01100_0110011;// and x12, x1, x2 -> x12 = x1(-100) & x2(3)
        */

        /*
        //rom[x] = 32'b imm7_ rs2 _rs1  _f3 _imm5 _op // S-Type
        rom[0] = 32'b0000000_00010_00000_000_00000_0100011;  // sb x2, 0(x0) 
        rom[1] = 32'b0000000_00010_00000_000_00101_0100011;  // sb x2, 5(x0) 
        rom[2] = 32'b0000000_00010_00000_010_01000_0100011;  // sw x2, 8(x0) 
        rom[3] = 32'b0000000_00010_00000_000_01010_0100011;  // sb x2, 10(x0)
        rom[4] = 32'b0000000_00010_00000_000_01111_0100011;  // sb x2, 15(x0)
        rom[5] = 32'b0000000_00010_00001_001_00101_0100011;  // sh x2, 5(x1)
        rom[6] = 32'b0000000_00010_00000_001_10110_0100011;  // sh x2, 22(x0)
        rom[7] = 32'b0000000_00010_00000_010_11000_0100011;  // sw x2, 24(x0)
        */

        /*
        //rom[x] = 32'b imm7_ rs2 _rs1  _f3 _imm5 _op // S-Type
        rom[0] = 32'b0000000_00001_00000_010_00000_0100011;  // sw x1, 0(x0)
        //rom[x] = 32'b imm12    _rs1  _f3 _rd   _op // L-Type
        rom[1] = 32'b000000000000_00000_010_00011_0000011;   // lw x3, 0(x0) 
        rom[2] = 32'b000000000000_00000_000_00100_0000011;   // lb x4, 0(x0) 
        rom[3] = 32'b000000000010_00000_000_00101_0000011;   // lb x5, 2(x0) 
        rom[4] = 32'b000000000010_00000_100_00110_0000011;   // lbu x6, 2(x0)
        rom[5] = 32'b000000000010_00000_001_00111_0000011;   // lh x7, 2(x0) 
        rom[6] = 32'b000000000010_00000_101_01000_0000011;   // lhu x8, 2(x0)
        */
        /*
        //rom[x] = 32'b imm       _rs1  _f3 _rd   _op   // I-Type
        rom[0] =  32'b000000001010_00001_000_00011_0010011;// addi x3, x1, 10 -> x3 = x1(-100) + x2(10)
        rom[1] =  32'b000000001010_00001_010_00100_0010011;// slti x4, x1, 10 -> x4 = x1(-100) < x2(10) ? 1 : 0
        rom[2] =  32'b000000001010_00001_011_00101_0010011;// sltiu x5, x1, 10 -> x5 = x1(-100) < x2(10) ? 1 : 0
        rom[3] =  32'b000000001010_00001_100_00110_0010011;// xori x6, x1, 10 -> x6 = x1(-100) ^ x2(10)
        rom[4] =  32'b000000001010_00001_110_00111_0010011;// ori x7, x1, 10 -> x7 = x1(-100) | x2(10)
        rom[5] =  32'b000000001010_00001_111_01000_0010011;// andi x8, x1, 10 -> x8 = x1(-100) & x2(10)
        rom[6] =  32'b0000000_00011_00001_001_01001_0010011;// slli x9, x1, 3 -> x9 = x1(-100) << x2(3)
        rom[7] =  32'b0000000_00011_00001_101_01010_0010011;// srli x10, x1, 3 -> x10 = x1(-100) >> x2(3)
        rom[8] =  32'b0100000_00011_00001_101_01011_0010011;// srai x11, x1, 3 -> x11 = x1(-100) >>> x2(3)
        */

        /*
        //rom[x] =  32'b imm7_ rs2 _rs1  _f3 _imm5 _op // B-Type
        //rom[x] = 32'b imm       _rs1  _f3 _rd   _op   // I-Type
        rom[0] =  32'b0000000_00010_00010_000_01000_1100011;// beq x2, x2, 8
        rom[1] =  32'b000000001010_00001_000_00011_0010011;//  addi x3, x1, 10 -> x3 = x1(-100) + 10
        rom[2] =  32'b0000000_00010_00010_001_01000_1100011;// bne x2, x2, 8
        rom[3] =  32'b000000001010_00001_010_00100_0010011;//  slti x4, x1, 10 -> x4 = x1(-100) < 10 ? 1 : 0
        rom[4] =  32'b0000000_00010_00001_100_01000_1100011;// blt x1, x2, 8
        rom[5] =  32'b000000001010_00001_011_00101_0010011;//  sltiu x5, x1, 10 -> x5 = x1(-100) < 10 ? 1 : 0
        rom[6] =  32'b0000000_00010_00001_101_01000_1100011;// bge x1, x2, 8
        rom[7] =  32'b000000001010_00001_100_00110_0010011;//  xori x6, x1, 10 -> x6 = x1(-100) ^ 10
        rom[8] =  32'b0000000_00010_00010_110_01000_1100011;// bltu x1, x2, 8
        rom[9] =  32'b000000001010_00001_110_00111_0010011;//  ori x7, x1, 10 -> x7 = x1(-100) | 10
        rom[10] =  32'b0000000_00010_00001_111_01000_1100011;//bgeu x1, x2, 8
        rom[11] =  32'b000000001010_00001_111_01000_0010011;// andi x8, x1, 10 -> x8 = x1(-100) & 10
        rom[12] =  32'b0000000_00011_00001_001_01001_0010011;//slli x9, x1, 3 -> x9 = x1(-100) << x2(3)
        */

        /*
        //rom[x] = 32'b imm       _rs1  _f3 _rd   _op   // I-Type
        rom[0] =  32'b000000000001_00001_000_00011_0010011; // addi x3, x1, 1
        rom[1] =  32'b0_0000000100_0_00000000_00100_1101111;// jal x4, 8
        rom[2] =  32'b000000000100_00010_111_00101_0010011; // andi x5, x2, 4
        rom[3] = 32'b000000000001_00010_110_00110_0010011;  // ori x6, x2, 1
        rom[4] = 32'b000000001100_00010_000_00111_1100111;  // jalr x7, x2, 24
        rom[5] = 32'b0000000_00010_00001_001_01000_0010011; // slli x8, x1, 2
        rom[6] = 32'b00000000000000000001_01001_0110111;    // lui  x9, 1 , 12
        rom[7] = 32'b00000000000000000001_01010_0010111;    // auipc x10 1, 12
        */

        /*
        
        //rom[x] = 32'b imm7_ rs2 _rs1  _f3 _imm5 _op // B-Type
        rom[5] = 32'b0000000_00010_00011_000_01100_1100011;  // beq x2, x3, 12
        //rom[x] = 32'b imm12    _rs1  _f3 _rd   _op // L-Type
        rom[6] = 32'b000000001000_00000_010_01000_0000011;  // lw x8, 8(x0)
        //rom[x] = 32'b imm12    _rs1  _f3 _rd   _op // I-Type
        rom[7] = 32'b000000000001_00001_000_01001_0010011;  // addi x9, x1, 1
        rom[8] = 32'b000000000100_00010_111_01010_0010011;  // andi x10, x2, 4
        rom[9] = 32'b000000000001_00010_110_01011_0010011;  // ori x11, x2, 1
        rom[10] = 32'b0000000_00010_00001_001_01100_0010011;  // slli x12, x1, 2
        */
    end
    assign data = rom[addr[31:2]];
endmodule